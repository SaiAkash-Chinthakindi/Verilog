`timescale 1ns / 1ps


module four_two_bit(A,y);
  input [3:0]A;
  output reg [1:0]y;
  
  always@(*)begin
    case(A)
      4'b1000 : y = 2'b11;
      4'b0100 : y = 2'b10;
      4'b0010 : y = 2'b01;
      4'b0001 : y = 2'b00;
      default : y = 2'b00;
    endcase
  end
  
endmodule
